module fadd(input logic [31:0] x1,
            input logic [31:0] x2,
            input logic clk,
            output logic [31:0] y
    );
    